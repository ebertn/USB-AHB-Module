mg69@ee215lnx10.ecn.purdue.edu.28936:1555451921