module tb_ahb_lite_slave ();



endmodule
