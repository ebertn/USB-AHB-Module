module state_controller (
	input wire clk,
	input wire nRst,
	
	input wire [6:0] haddr,
	input wire [1:0] htrans,
	input wire [1:0] hsize,
	input wire hwrite,
	input wire hsel,
	
	output reg [1:0] state,
	output reg storeTxData,
	output reg getRxData,
	output reg hresp,
	output reg hready,
	output wire [1:0] dataSize,
	output logic txPacketSizeChanged
);

// localparams
localparam IDLE = 2'b00;
localparam WRITE = 2'b01;
localparam READ = 2'b10;
localparam ERROR = 2'b11;

// internal signals
reg [1:0] nextState;

// Small Assignments
assign dataSize = hsize;
assign hresp = ((state == ERROR) || (nextState == ERROR)) ? 1'b1 : 1'b0;
assign hready = (nextState == ERROR) ? 1'b0 : 1'b1;

// Next State Logic
always_comb begin
	storeTxData = 1'b0;
	getRxData = 1'b0;
	nextState = IDLE;
	txPacketSizeChanged = 1'b0;

	if (hsel && (htrans != IDLE)) begin
		if (hsize == 2'b11) begin
			nextState = ERROR;
			
		end else if (hwrite) begin
			if ((haddr >= 7'h00) && (haddr < 7'h40)) begin
				storeTxData = 1'b1;
				nextState = WRITE;
			end else if ((haddr == 7'h48) && (hsize == 2'b00)) begin
				nextState = WRITE;
				txPacketSizeChanged = 1'b1;
			end else begin
				nextState = ERROR;
			end
			
		end else if (!hwrite) begin
			if ((haddr >= 7'h00) && (haddr < 7'h40)) begin
				getRxData = 1'b1;
				nextState = READ;
			end else if (((haddr == 7'h40) || (haddr == 7'h41)) && ((hsize == 2'b01) || (hsize == 2'b00))) begin
				nextState = READ;
			end else if (((haddr == 7'h42) || (haddr == 7'h43)) && ((hsize == 2'b01) || (hsize == 2'b00))) begin
				nextState = READ;
			end else if (((haddr == 7'h44) || (haddr == 7'h48)) && (hsize == 2'b00)) begin
				nextState = READ;
			end else begin
				nextState = ERROR;
			end
			
		end else begin
			nextState = ERROR;
		end
	end
end

// Register for State
always_ff @(posedge clk, negedge nRst) begin
	if (nRst == 1'b0) begin
		state <= IDLE;
	end else begin
		state <= nextState;
	end
end

endmodule
